package htfft{{suffix}}_params is
  constant INPUT_WIDTH: positive := {{input_width}};
  constant OUTPUT_WIDTH: positive := {{output_width}};
  constant N: positive := {{n}};
  constant SPCC: positive := {{spcc}};

end package;
